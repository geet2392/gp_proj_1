Welcome to project modified just now:w
