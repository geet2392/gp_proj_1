Welcome to project
added line at diffrent pos
line 3 added 


