Welcome to project
added line at diffrent pos
line 3 added 


<<<<<<< HEAD
line 5 added


=======
>>>>>>> f7458b65327b66154e3f0abaa882c087a5c8e350
