Welcome to project
added line at diffrent pos
