Welcome to project
added line at diffrent pos
line 3 added 


line 5 added


